   REGISTER_EN        = 1         ,
   REGISTER_EPDATA    = 0         ,
   PKTCNTWD           = 9        ,
   ADDR_SIZE          = 32        ,
   DATA_SIZE          = 32        ,
  START_EPT_HADDR    = 32'h00_0920 ,
   END_EPT_HADDR      = 32'h00_0D9C ,
   START_REG_HADDR1   = 32'h00_0800 ,  
   END_REG_HADDR1     = 32'h00_091B 
