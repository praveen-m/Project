   ADDR_SIZE          = 32        ,
   DATA_SIZE          = 32        , 
   REGISTER_EN        = 1         ,
   REGISTER_EPDATA    = 0         ,
   PKTCNTWD           = 9         ,
   BYPASS             = 1           ,
   START_EPT_HADDR    = 32'h00_0920 ,
   END_EPT_HADDR      = 32'h00_0D9C ,
   START_REG_HADDR1   = 32'h00_0800 ,  
   END_REG_HADDR1     = 32'h00_091B , 
   //register address parameter
   SUSP_CTRL          = 32'h0800  ,
   RESET_CTRL         = 32'h0804  ,
   DEV_CTRL1          = 32'h0808  ,
   DEV_CTRL2          = 32'h080C  ,
   DEV_STAT1          = 32'h0810  ,
   DEV_STAT2          = 32'h0814  ,
   CTRL_EP_CMD_REG    = 32'h0820  ,
   CTRL_EP_RD_ADDR    = 32'h0824  ,
   MEM_SEG_ADDR       = 32'h082C  ,
   DMA_TX_ADDR        = 32'h0830  ,
   EP_WR_ADDR         = 32'h0834  ,
   EBUF_TX_CTRL1      = 32'h0838  ,
   EBUF_TX_CTRL2      = 32'h083C  ,
   DMA_RX_ADDR        = 32'h0840  ,
   EBUF_RX_CTRL1      = 32'h0844  ,
   EBUF_RX_CTRL2      = 32'h0848  ,
   SOF_COUNT          = 32'h0850  ,
   SOF_CTRL           = 32'h0854  ,
   SOF_TIMER_SET      = 32'h0858  ,
   SETUP_CMD1         = 32'h0860  ,
   SETUP_CMD2         = 32'h0864  ,
   TIMER_CTRL1        = 32'h0870  ,
   TIMER_CTRL2        = 32'h0874  ,
   TIMER_CTRL3        = 32'h0878  ,
   TIMER_CTRL4        = 32'h087C  ,
   TIMER_CTRL5        = 32'h0880  ,
   TIMER_CTRL6        = 32'h0884  ,
   TIMER_CTRL7        = 32'h0888  ,
   TIMER_CTRL8        = 32'h088C  ,
   TIMER_CTRL9        = 32'h0890  ,
   TIMER_CTRL10       = 32'h0894  ,
   TIMER_CTRL11       = 32'h0898  ,
   TIMER_CTRL12       = 32'h089C  ,
   TIMER_CTRL13       = 32'h08A0  ,
   TIMER_CTRL14       = 32'h08A4  ,
   TIMER_CTRL15       = 32'h08A8  ,
   TIMER_CTRL16       = 32'h08AC  ,
   TIMER_CTRL17       = 32'h08B0  ,
   TIMER_CTRL18       = 32'h08B4  ,
   TIMER_CTRL19       = 32'h08B8  ,
   TIMER_CTRL20       = 32'h08BC  ,
   INTR_MASK_PRI      = 32'h08C0  ,
   INTR_MASK_SEC      = 32'h08C8  ,
   INTR_STATUS_PRI    = 32'h08D0  ,
   INTR_STATUS_SEC    = 32'h08D8  ,
   INTR_DATA1_PRI     = 32'h08E0  ,
   INTR_DATA2_PRI     = 32'h08E4  ,
   INTR_DATA1_SEC     = 32'h08EC  ,
   INTR_DATA2_SEC     = 32'h08F0  ,
   TEST_CTRL          = 32'h08F8  ,
   USB_TRANS_CTRL     = 32'h0900  ,
   USB_TX_TRANS_DATA1 = 32'h0904  ,
   USB_TX_TRANS_DATA2 = 32'h0908  ,
   USB_TX_TRANS_DATA3 = 32'h090C  ,
   USB_RX_TRANS_DATA1 = 32'h0910  ,
   USB_RX_TRANS_DATA2 = 32'h0914  ,
   USB_RX_TRANS_DATA3 = 32'h0918  ,
   // endpoint data address parameter
   EPT0_SA           =  32'h0920  ,
   EPT0_EA           =  32'h0924  ,
   EPT0_CR1          =  32'h0928  ,
   EPT0_CR2          =  32'h092C  ,
   EPT0_WPTR         =  32'h0930  ,
   EPT0_RPTR         =  32'h0934  ,
   EPT0_STAT         =  32'h093C  ,
   EPT1_SA           =  32'h0940  ,
   EPT1_EA           =  32'h0944  ,
   EPT1_CR1          =  32'h0948  ,
   EPT1_CR2          =  32'h094C  ,
   EPT1_WPTR         =  32'h0950  ,
   EPT1_RPTR         =  32'h0954  ,
   EPT1_STAT         =  32'h095C  ,
   EPT2_SA           =  32'h0960  ,
   EPT2_EA           =  32'h0964  ,
   EPT2_CR1          =  32'h0968  ,
   EPT2_CR2          =  32'h096C  ,
   EPT2_WPTR         =  32'h0970  ,
   EPT2_RPTR         =  32'h0974  ,
   EPT2_STAT         =  32'h097C  ,
   EPT3_SA           =  32'h0980  ,
   EPT3_EA           =  32'h0984  ,
   EPT3_CR1          =  32'h0988  ,
   EPT3_CR2          =  32'h098C  ,
   EPT3_WPTR         =  32'h0990  ,
   EPT3_RPTR         =  32'h0994  ,
   EPT3_STAT         =  32'h099C  ,
   EPT4_SA           =  32'h09A0  ,
   EPT4_EA           =  32'h09A4  ,
   EPT4_CR1          =  32'h09A8  ,
   EPT4_CR2          =  32'h09AC  ,
   EPT4_WPTR         =  32'h09B0  ,
   EPT4_RPTR         =  32'h09B4  ,
   EPT4_STAT         =  32'h09BC  ,
   EPT5_SA           =  32'h09C0  ,
   EPT5_EA           =  32'h09C4  ,
   EPT5_CR1          =  32'h09C8  ,
   EPT5_CR2          =  32'h09CC  ,
   EPT5_WPTR         =  32'h09D0  ,
   EPT5_RPTR         =  32'h09D4  ,
   EPT5_STAT         =  32'h09DC  ,
   EPT6_SA           =  32'h09E0  ,
   EPT6_EA           =  32'h09E4  ,
   EPT6_CR1          =  32'h09E8  ,
   EPT6_CR2          =  32'h09EC  ,
   EPT6_WPTR         =  32'h09F0  ,
   EPT6_RPTR         =  32'h09F4  ,
   EPT6_STAT         =  32'h09FC  ,
   EPT7_SA           =  32'h0A00  ,
   EPT7_EA           =  32'h0A04  ,
   EPT7_CR1          =  32'h0A08  ,
   EPT7_CR2          =  32'h0A0C  ,
   EPT7_WPTR         =  32'h0A10  ,
   EPT7_RPTR         =  32'h0A14  ,
   EPT7_STAT         =  32'h0A1C  ,
   EPT8_SA           =  32'h0A20  ,
   EPT8_EA           =  32'h0A24  ,
   EPT8_CR1          =  32'h0A28  ,
   EPT8_CR2          =  32'h0A2C  ,
   EPT8_WPTR         =  32'h0A30  ,
   EPT8_RPTR         =  32'h0A34  ,
   EPT8_STAT         =  32'h0A3C  ,
   EPT9_SA           =  32'h0A40  ,
   EPT9_EA           =  32'h0A44  ,
   EPT9_CR1          =  32'h0A48  ,
   EPT9_CR2          =  32'h0A4C  ,
   EPT9_WPTR         =  32'h0A50  ,
   EPT9_RPTR         =  32'h0A54  ,
   EPT9_STAT         =  32'h0A5C  ,
   EPT10_SA          =  32'h0A60  ,
   EPT10_EA          =  32'h0A64  ,
   EPT10_CR1         =  32'h0A68  ,
   EPT10_CR2         =  32'h0A6C  ,
   EPT10_WPTR        =  32'h0A70  ,
   EPT10_RPTR        =  32'h0A74  ,
   EPT10_STAT        =  32'h0A7C  ,
   EPT11_SA          =  32'h0A80  ,
   EPT11_EA          =  32'h0A84  ,
   EPT11_CR1         =  32'h0A88  ,
   EPT11_CR2         =  32'h0A8C  ,
   EPT11_WPTR        =  32'h0A90  ,
   EPT11_RPTR        =  32'h0A94  ,
   EPT11_STAT        =  32'h0A9C  ,
   EPT12_SA          =  32'h0AA0  ,
   EPT12_EA          =  32'h0AA4  ,
   EPT12_CR1         =  32'h0AA8  ,
   EPT12_CR2         =  32'h0AAC  ,
   EPT12_WPTR        =  32'h0AB0  ,
   EPT12_RPTR        =  32'h0AB4  ,
   EPT12_STAT        =  32'h0ABC  ,
   EPT13_SA          =  32'h0AC0  ,
   EPT13_EA          =  32'h0AC4  ,
   EPT13_CR1         =  32'h0AC8  ,
   EPT13_CR2         =  32'h0ACC  ,
   EPT13_WPTR        =  32'h0AD0  ,
   EPT13_RPTR        =  32'h0AD4  ,
   EPT13_STAT        =  32'h0ADC  ,
   EPT14_SA          =  32'h0AE0  ,
   EPT14_EA          =  32'h0AE4  ,
   EPT14_CR1         =  32'h0AE8  ,
   EPT14_CR2         =  32'h0AEC  ,
   EPT14_WPTR        =  32'h0AF0  ,
   EPT14_RPTR        =  32'h0AF4  ,
   EPT14_STAT        =  32'h0AFC  ,
   EPT15_SA          =  32'h0B00  ,
   EPT15_EA          =  32'h0B04  ,
   EPT15_CR1         =  32'h0B08  ,
   EPT15_CR2         =  32'h0B0C  ,
   EPT15_WPTR        =  32'h0B10  ,
   EPT15_RPTR        =  32'h0B14  ,
   EPT15_STAT        =  32'h0B1C  ,
   EPT16_SA          =  32'h0B20  ,
   EPT16_EA          =  32'h0B24  ,
   EPT16_CR1         =  32'h0B28  ,
   EPT16_CR2         =  32'h0B2C  ,
   EPT16_WPTR        =  32'h0B30  ,
   EPT16_RPTR        =  32'h0B34  ,
   EPT16_ARPTR       =  32'h0B38  ,
   EPT16_STAT        =  32'h0B3C  ,
   EPT17_SA          =  32'h0B40  ,
   EPT17_EA          =  32'h0B44  ,
   EPT17_CR1         =  32'h0B48  ,
   EPT17_CR2         =  32'h0B4C  ,
   EPT17_WPTR        =  32'h0B50  ,
   EPT17_RPTR        =  32'h0B54  ,
   EPT17_ARPTR       =  32'h0B58  ,
   EPT17_STAT        =  32'h0B5C  ,
   EPT18_SA          =  32'h0B60  ,
   EPT18_EA          =  32'h0B64  ,
   EPT18_CR1         =  32'h0B68  ,
   EPT18_CR2         =  32'h0B6C  ,
   EPT18_WPTR        =  32'h0B70  ,
   EPT18_RPTR        =  32'h0B74  ,
   EPT18_ARPTR       =  32'h0B78  ,
   EPT18_STAT        =  32'h0B7C  ,
   EPT19_SA          =  32'h0B80  ,
   EPT19_EA          =  32'h0B84  ,
   EPT19_CR1         =  32'h0B88  ,
   EPT19_CR2         =  32'h0B8C  ,
   EPT19_WPTR        =  32'h0B90  ,
   EPT19_RPTR        =  32'h0B94  ,
   EPT19_ARPTR       =  32'h0B98  ,
   EPT19_STAT        =  32'h0B9C  ,
   EPT20_SA          =  32'h0BA0  ,
   EPT20_EA          =  32'h0BA4  ,
   EPT20_CR1         =  32'h0BA8  ,
   EPT20_CR2         =  32'h0BAC  ,
   EPT20_WPTR        =  32'h0BB0  ,
   EPT20_RPTR        =  32'h0BB4  ,
   EPT20_ARPTR       =  32'h0BB8  ,
   EPT20_STAT        =  32'h0BBC  ,
   EPT21_SA          =  32'h0BC0  ,
   EPT21_EA          =  32'h0BC4  ,
   EPT21_CR1         =  32'h0BC8  ,
   EPT21_CR2         =  32'h0BCC  ,
   EPT21_WPTR        =  32'h0BD0  ,
   EPT21_RPTR        =  32'h0BD4  ,
   EPT21_ARPTR       =  32'h0BD8  ,
   EPT21_STAT        =  32'h0BDC  ,
   EPT22_SA          =  32'h0BE0  ,
   EPT22_EA          =  32'h0BE4  ,
   EPT22_CR1         =  32'h0BE8  ,
   EPT22_CR2         =  32'h0BEC  ,
   EPT22_WPTR        =  32'h0BF0  ,
   EPT22_RPTR        =  32'h0BF4  ,
   EPT22_ARPTR       =  32'h0BF8  ,
   EPT22_STAT        =  32'h0BFC  ,
   EPT23_SA          =  32'h0C00  ,
   EPT23_EA          =  32'h0C04  ,
   EPT23_CR1         =  32'h0C08  ,
   EPT23_CR2         =  32'h0C0C  ,
   EPT23_WPTR        =  32'h0C10  ,
   EPT23_RPTR        =  32'h0C14  ,
   EPT23_ARPTR       =  32'h0C18  ,
   EPT23_STAT        =  32'h0C1C  ,
   EPT24_SA          =  32'h0C20  ,
   EPT24_EA          =  32'h0C24  ,
   EPT24_CR1         =  32'h0C28  ,
   EPT24_CR2         =  32'h0C2C  ,
   EPT24_WPTR        =  32'h0C30  ,
   EPT24_RPTR        =  32'h0C34  ,
   EPT24_ARPTR       =  32'h0C38  ,
   EPT24_STAT        =  32'h0C3C  ,
   EPT25_SA          =  32'h0C40  ,
   EPT25_EA          =  32'h0C44  ,
   EPT25_CR1         =  32'h0C48  ,
   EPT25_CR2         =  32'h0C4C  ,
   EPT25_WPTR        =  32'h0C50  ,
   EPT25_RPTR        =  32'h0C54  ,
   EPT25_ARPTR       =  32'h0C58  ,
   EPT25_STAT        =  32'h0C5C  ,
   EPT26_SA          =  32'h0C60  ,
   EPT26_EA          =  32'h0C64  ,
   EPT26_CR1         =  32'h0C68  ,
   EPT26_CR2         =  32'h0C6C  ,
   EPT26_WPTR        =  32'h0C70  ,
   EPT26_RPTR        =  32'h0C74  ,
   EPT26_ARPTR       =  32'h0C78  ,
   EPT26_STAT        =  32'h0C7C  ,
   EPT27_SA          =  32'h0C80  ,
   EPT27_EA          =  32'h0C84  ,
   EPT27_CR1         =  32'h0C88  ,
   EPT27_CR2         =  32'h0C8C  ,
   EPT27_WPTR        =  32'h0C90  ,
   EPT27_RPTR        =  32'h0C94  ,
   EPT27_ARPTR       =  32'h0C98  ,
   EPT27_STAT        =  32'h0C9C  ,
   EPT28_SA          =  32'h0CA0  ,
   EPT28_EA          =  32'h0CA4  ,
   EPT28_CR1         =  32'h0CA8  ,
   EPT28_CR2         =  32'h0CAC  ,
   EPT28_WPTR        =  32'h0CB0  ,
   EPT28_RPTR        =  32'h0CB4  ,
   EPT28_ARPTR       =  32'h0CB8  ,
   EPT28_STAT        =  32'h0CBC  ,
   EPT29_SA          =  32'h0CC0  ,
   EPT29_EA          =  32'h0CC4  ,
   EPT29_CR1         =  32'h0CC8  ,
   EPT29_CR2         =  32'h0CCC  ,
   EPT29_WPTR        =  32'h0CD0  ,
   EPT29_RPTR        =  32'h0CD4  ,
   EPT29_ARPTR       =  32'h0CD8  ,
   EPT29_STAT        =  32'h0CDC  ,
   EPT30_SA          =  32'h0CE0  ,
   EPT30_EA          =  32'h0CE4  ,
   EPT30_CR1         =  32'h0CE8  ,
   EPT30_CR2         =  32'h0CEC  ,
   EPT30_WPTR        =  32'h0CF0  ,
   EPT30_RPTR        =  32'h0CF4  ,
   EPT30_ARPTR       =  32'h0CF8  ,
   EPT30_STAT        =  32'h0CFC  ,
   EPT31_SA          =  32'h0D00  ,
   EPT31_EA          =  32'h0D04  ,
   EPT31_CR1         =  32'h0D08  ,
   EPT31_CR2         =  32'h0D0C  ,
   EPT31_WPTR        =  32'h0D10  ,
   EPT31_RPTR        =  32'h0D14  ,
   EPT31_ARPTR       =  32'h0D18  ,
   EPT31_STAT        =  32'h0D1C  ,
   EPT0_FULLBUFCNT   =  32'h0D20  ,
   EPT1_FULLBUFCNT   =  32'h0D24  ,
   EPT2_FULLBUFCNT   =  32'h0D28  ,
   EPT3_FULLBUFCNT   =  32'h0D2C  ,
   EPT4_FULLBUFCNT   =  32'h0D30  ,
   EPT5_FULLBUFCNT   =  32'h0D34  ,
   EPT6_FULLBUFCNT   =  32'h0D38  ,
   EPT7_FULLBUFCNT   =  32'h0D3C  ,
   EPT8_FULLBUFCNT   =  32'h0D40  ,
   EPT9_FULLBUFCNT   =  32'h0D44  ,
   EPT10_FULLBUFCNT  =  32'h0D48  ,
   EPT11_FULLBUFCNT  =  32'h0D4C  ,
   EPT12_FULLBUFCNT  =  32'h0D50  ,
   EPT13_FULLBUFCNT  =  32'h0D54  ,
   EPT14_FULLBUFCNT  =  32'h0D58  ,
   EPT15_FULLBUFCNT  =  32'h0D5C  ,
   EPT16_FULLBUFCNT  =  32'h0D60  ,
   EPT17_FULLBUFCNT  =  32'h0D64  ,
   EPT18_FULLBUFCNT  =  32'h0D68  ,
   EPT19_FULLBUFCNT  =  32'h0D6C  ,
   EPT20_FULLBUFCNT  =  32'h0D70  ,
   EPT21_FULLBUFCNT  =  32'h0D74  ,
   EPT22_FULLBUFCNT  =  32'h0D78  ,
   EPT23_FULLBUFCNT  =  32'h0D7C  ,
   EPT24_FULLBUFCNT  =  32'h0D80  ,
   EPT25_FULLBUFCNT  =  32'h0D84  ,
   EPT26_FULLBUFCNT  =  32'h0D88  ,
   EPT27_FULLBUFCNT  =  32'h0D8C  ,
   EPT28_FULLBUFCNT  =  32'h0D90  ,
   EPT29_FULLBUFCNT  =  32'h0D94  ,
   EPT30_FULLBUFCNT  =  32'h0D98  ,
   EPT31_FULLBUFCNT  =  32'h0D9C  
                             
